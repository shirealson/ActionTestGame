LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.MATH_REAL.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY button_scan IS
PORT(
      game_clk:IN STD_LOGIC;
	  kbrow:IN STD_LOGIC_VECTOR(3 downto 0);
	  button_output : out std_logic_vector(3 downto 0)
);
END ENTITY button_scan;

architecture a of button_scan is
	SIGNAL up,down,left,right : std_logic:='0';
	SIGNAL kbcols:STD_LOGIC_VECTOR(0 TO 3); 
	
	
begin	

	process(game_clk)
	begin
		if game_clk'event and game_clk = '1' then
			if kbrow = "0111" then
				up <= '1'; 
			else 
				up <= '0';
			end if;
			
			if kbrow = "1011" then
				left <= '1'; 
			else 
				left <= '0';
			end if;
			
			if kbrow = "1101" then
				right <= '1'; 
			else 
				right <= '0';
			end if;
			
			if kbrow = "1110" then
				down <= '1'; 
			else 
				down <= '0';
			end if;
		end if;
	end process;
	--------------------------------------------------------------------------------------------------------------
--�������������
	OUTPUT_KEY : process(up,down,left,right)
	begin
	if up = '1' then
		button_output <= "1000";
	elsif down = '1' then
		button_output <= "0100";
	elsif left = '1' then
		button_output <= "0010";
	elsif right = '1' then
		button_output <= "0001";
	else
		button_output <= "0000";
	end if;
	end process OUTPUT_KEY; 


end a;
	
	
